module hello;
    initial $display ("Hello world!");
endmodule
